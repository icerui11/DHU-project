----------------------------------------------------------------------------------------------------------------------------------
-- File Description  --
----------------------------------------------------------------------------------------------------------------------------------
-- @ File Name				:	router_oneShyloc_top.vhd
-- @ Engineer				:	Rui Yin
-- @ Role					:	FPGA Engineer
-- @ Company				:	4Links ltd
-- @ Date					: 	12/12/2024

-- @ VHDL Version			:   1987, 1993, 2008
-- @ Supported Toolchain	:	libero
-- @ Target Device			: 	SmartFusion2

-- @ Revision #				:	1

-- File Description         :

-- Document Number			:  xxx-xxxx-xxx
----------------------------------------------------------------------------------------------------------------------------------
-- Library Declarations  --
----------------------------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

----------------------------------------------------------------------------------------------------------------------------------
-- Package Declarations --
----------------------------------------------------------------------------------------------------------------------------------
context work.router_context;

----------------------------------------------------------------------------------------------------------------------------------
-- Entity Declarations --
----------------------------------------------------------------------------------------------------------------------------------
entity router_oneShyloc_top is
    generic(
		g_clock_freq	: real 					:= c_spw_clk_freq;
        g_num_ports 	: natural range 1 to 32 := c_num_ports;
		g_mode			: string				:= c_port_mode;
		g_is_fifo		: t_dword 				:= c_fifo_ports;
		g_priority		: string 				:= c_priority;
		g_ram_style 	: string				:= c_ram_style 
    );
	port( 
		clk_in		    : in 	std_logic := '0';		-- router clock input 
		rst_in			: in 	std_logic := '0';		-- reset input, active high

		Din_p  			: in 	std_logic_vector(1 to g_num_ports-1)	:= (others => '0');
		Sin_p           : in 	std_logic_vector(1 to g_num_ports-1)	:= (others => '0');
		Dout_p          : out 	std_logic_vector(1 to g_num_ports-1)	:= (others => '0');
		Sout_p          : out 	std_logic_vector(1 to g_num_ports-1)	:= (others => '0');

		--port_connected	: out 	std_logic_vector(31 downto 1) := (others => '0');	-- High when "connected" May want to map these to LEDs
		
		spw_en_pinout	: out	std_logic_vector(1 to g_num_ports-1) := (others => '0')

    );
end router_oneShyloc_top;


---------------------------------------------------------------------------------------------------------------------------------
-- Code Description & Developer Notes --
---------------------------------------------------------------------------------------------------------------------------------


architecture rtl of router_oneShyloc_top is

	----------------------------------------------------------------------------------------------------------------------------
	-- Constant Declarations --
	----------------------------------------------------------------------------------------------------------------------------

	----------------------------------------------------------------------------------------------------------------------------
	-- Type Declarations --
	----------------------------------------------------------------------------------------------------------------------------
	
	----------------------------------------------------------------------------------------------------------------------------
	-- Function Declarations --
	----------------------------------------------------------------------------------------------------------------------------

	----------------------------------------------------------------------------------------------------------------------------
	-- Entity Declarations --
	----------------------------------------------------------------------------------------------------------------------------
	
	----------------------------------------------------------------------------------------------------------------------------
	-- Component Declarations --
	----------------------------------------------------------------------------------------------------------------------------
	
	----------------------------------------------------------------------------------------------------------------------------
	-- Signal Declarations --
	----------------------------------------------------------------------------------------------------------------------------
    
	----------------------------------------------------------------------------------------------------------------------------
	-- Variable Declarations --
	----------------------------------------------------------------------------------------------------------------------------

	----------------------------------------------------------------------------------------------------------------------------
	-- Alias Declarations --
	----------------------------------------------------------------------------------------------------------------------------
	
	----------------------------------------------------------------------------------------------------------------------------
	-- Attribute Declarations --
	----------------------------------------------------------------------------------------------------------------------------
	
begin
	
	----------------------------------------------------------------------------------------------------------------------------
	-- Entity Instantiations --
	----------------------------------------------------------------------------------------------------------------------------
	router_inst: entity work.router_top_level_RTG4(rtl)	-- instantiate SpaceWire Router 
	generic map(
		g_clock_freq 	=> g_clock_freq,
		g_num_ports 	=> g_num_ports,
		g_is_fifo 		=> g_is_fifo,
		g_mode			=> "single",					-- custom mode, we're instantiating SpaceWire in this top-level architecture
		g_priority 		=> g_priority,
		g_ram_style 	=> g_ram_style
	)
	port map( 

		router_clk              => clk_in,
		rst_in					=> rst_in,	 
	
		DDR_din_r				=> '0',	
		DDR_din_f   			=> '0',  
		DDR_sin_r   			=> '0',  
		DDR_sin_f   			=> '0',  
		SDR_Dout				=> open,
		SDR_Sout				=> open,
		
		Din_p               	=> Din_p, 
		Din_n               	=> '0', 
		Sin_p               	=> Sin_p, 
		Sin_n               	=> '0', 
		Dout_p              	=> Dout_p, 
		Dout_n              	=> open, 
		Sout_p              	=> Sout_p, 
		Sout_n              	=> open,  

		spw_fifo_in             => spw_fifo_in,
		spw_fifo_out	        => spw_fifo_out,
		
		Port_Connected			=> open
	);

    
	----------------------------------------------------------------------------------------------------------------------------
	-- Component Instantiations --
	----------------------------------------------------------------------------------------------------------------------------

	----------------------------------------------------------------------------------------------------------------------------
	-- Asynchronous Signal Assignments --
	----------------------------------------------------------------------------------------------------------------------------

	----------------------------------------------------------------------------------------------------------------------------
	-- Synchronous Processes --
	----------------------------------------------------------------------------------------------------------------------------
end rtl;