--============================================================================--
-- Design unit  : rom_data
--
-- File name    : allones_h8w7b5_8int_le.bip.vhd
--
-- Purpose      : data for the ROM
--
-- Note         :
--
-- Library      : shyloc_utils
--
-- Author       : Rui Yin
--
-- Instantiates : 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

package ROM_Package is
	
    constant width	: integer := 8;
    constant depth : integer:= 3072;
    constant addr : integer := 10;
    type ROM_ARRAY is array (0 to depth-1) of STD_LOGIC_VECTOR(width-1 downto 0);
    constant ROM_CONTENT: ROM_ARRAY := (
    0 => X"00",
    1 => X"01",
    2 => X"02",
    3 => X"03",
    4 => X"04",
    5 => X"05",
    6 => X"06",
    7 => X"07",
    8 => X"08",
    9 => X"09",
    10 => X"0A",
    11 => X"0B",
    12 => X"0C",
    13 => X"0D",
    14 => X"0E",
    15 => X"0F",
    16 => X"10",
    17 => X"11",
    18 => X"12",
    19 => X"13",
    20 => X"14",
    21 => X"15",
    22 => X"16",
    23 => X"17",
    24 => X"18",
    25 => X"19",
    26 => X"1A",
    27 => X"1B",
    28 => X"1C",
    29 => X"1D",
    30 => X"1E",
    31 => X"1F",
    32 => X"20",
    33 => X"21",
    34 => X"22",
    35 => X"23",
    36 => X"24",
    37 => X"25",
    38 => X"26",
    39 => X"27",
    40 => X"28",
    41 => X"29",
    42 => X"2A",
    43 => X"2B",
    44 => X"2C",
    45 => X"2D",
    46 => X"2E",
    47 => X"2F",
    48 => X"30",
    49 => X"31",
    50 => X"32",
    51 => X"33",
    52 => X"34",
    53 => X"35",
    54 => X"36",
    55 => X"37",
    56 => X"38",
    57 => X"39",
    58 => X"3A",
    59 => X"3B",
    60 => X"3C",
    61 => X"3D",
    62 => X"3E",
    63 => X"3F",
    64 => X"40",
    65 => X"41",
    66 => X"42",
    67 => X"43",
    68 => X"44",
    69 => X"45",
    70 => X"46",
    71 => X"47",
    72 => X"48",
    73 => X"49",
    74 => X"4A",
    75 => X"4B",
    76 => X"4C",
    77 => X"4D",
    78 => X"4E",
    79 => X"4F",
    80 => X"50",
    81 => X"51",
    82 => X"52",
    83 => X"53",
    84 => X"54",
    85 => X"55",
    86 => X"56",
    87 => X"57",
    88 => X"58",
    89 => X"59",
    90 => X"5A",
    91 => X"5B",
    92 => X"5C",
    93 => X"5D",
    94 => X"5E",
    95 => X"5F",
    96 => X"60",
    97 => X"61",
    98 => X"62",
    99 => X"63",
    100 => X"64",
    101 => X"65",
    102 => X"66",
    103 => X"67",
    104 => X"68",
    105 => X"69",
    106 => X"6A",
    107 => X"6B",
    108 => X"6C",
    109 => X"6D",
    110 => X"6E",
    111 => X"6F",
    112 => X"70",
    113 => X"71",
    114 => X"72",
    115 => X"73",
    116 => X"74",
    117 => X"75",
    118 => X"76",
    119 => X"77",
    120 => X"78",
    121 => X"79",
    122 => X"7A",
    123 => X"7B",
    124 => X"7C",
    125 => X"7D",
    126 => X"7E",
    127 => X"7F",
    128 => X"80",
    129 => X"81",
    130 => X"82",
    131 => X"83",
    132 => X"84",
    133 => X"85",
    134 => X"86",
    135 => X"87",
    136 => X"88",
    137 => X"89",
    138 => X"8A",
    139 => X"8B",
    140 => X"8C",
    141 => X"8D",
    142 => X"8E",
    143 => X"8F",
    144 => X"90",
    145 => X"91",
    146 => X"92",
    147 => X"93",
    148 => X"94",
    149 => X"95",
    150 => X"96",
    151 => X"97",
    152 => X"98",
    153 => X"99",
    154 => X"9A",
    155 => X"9B",
    156 => X"9C",
    157 => X"9D",
    158 => X"9E",
    159 => X"9F",
    160 => X"A0",
    161 => X"A1",
    162 => X"A2",
    163 => X"A3",
    164 => X"A4",
    165 => X"A5",
    166 => X"A6",
    167 => X"A7",
    168 => X"A8",
    169 => X"A9",
    170 => X"AA",
    171 => X"AB",
    172 => X"AC",
    173 => X"AD",
    174 => X"AE",
    175 => X"AF",
    176 => X"B0",
    177 => X"B1",
    178 => X"B2",
    179 => X"B3",
    180 => X"B4",
    181 => X"B5",
    182 => X"B6",
    183 => X"B7",
    184 => X"B8",
    185 => X"B9",
    186 => X"BA",
    187 => X"BB",
    188 => X"BC",
    189 => X"BD",
    190 => X"BE",
    191 => X"BF",
    192 => X"C0",
    193 => X"C1",
    194 => X"C2",
    195 => X"C3",
    196 => X"C4",
    197 => X"C5",
    198 => X"C6",
    199 => X"C7",
    200 => X"C8",
    201 => X"C9",
    202 => X"CA",
    203 => X"CB",
    204 => X"CC",
    205 => X"CD",
    206 => X"CE",
    207 => X"CF",
    208 => X"D0",
    209 => X"D1",
    210 => X"D2",
    211 => X"D3",
    212 => X"D4",
    213 => X"D5",
    214 => X"D6",
    215 => X"D7",
    216 => X"D8",
    217 => X"D9",
    218 => X"DA",
    219 => X"DB",
    220 => X"DC",
    221 => X"DD",
    222 => X"DE",
    223 => X"DF",
    224 => X"E0",
    225 => X"E1",
    226 => X"E2",
    227 => X"E3",
    228 => X"E4",
    229 => X"E5",
    230 => X"E6",
    231 => X"E7",
    232 => X"E8",
    233 => X"E9",
    234 => X"EA",
    235 => X"EB",
    236 => X"EC",
    237 => X"ED",
    238 => X"EE",
    239 => X"EF",
    240 => X"F0",
    241 => X"F1",
    242 => X"F2",
    243 => X"F3",
    244 => X"F4",
    245 => X"F5",
    246 => X"F6",
    247 => X"F7",
    248 => X"F8",
    249 => X"F9",
    250 => X"FA",
    251 => X"FB",
    252 => X"FC",
    253 => X"FD",
    254 => X"FE",
    255 => X"FF",
    256 => X"00",
    257 => X"01",
    258 => X"02",
    259 => X"03",
    260 => X"04",
    261 => X"05",
    262 => X"06",
    263 => X"07",
    264 => X"08",
    265 => X"09",
    266 => X"0A",
    267 => X"0B",
    268 => X"0C",
    269 => X"0D",
    270 => X"0E",
    271 => X"0F",
    272 => X"10",
    273 => X"11",
    274 => X"12",
    275 => X"13",
    276 => X"14",
    277 => X"15",
    278 => X"16",
    279 => X"17",
    280 => X"18",
    281 => X"19",
    282 => X"1A",
    283 => X"1B",
    284 => X"1C",
    285 => X"1D",
    286 => X"1E",
    287 => X"1F",
    288 => X"20",
    289 => X"21",
    290 => X"22",
    291 => X"23",
    292 => X"24",
    293 => X"25",
    294 => X"26",
    295 => X"27",
    296 => X"28",
    297 => X"29",
    298 => X"2A",
    299 => X"2B",
    300 => X"2C",
    301 => X"2D",
    302 => X"2E",
    303 => X"2F",
    304 => X"30",
    305 => X"31",
    306 => X"32",
    307 => X"33",
    308 => X"34",
    309 => X"35",
    310 => X"36",
    311 => X"37",
    312 => X"38",
    313 => X"39",
    314 => X"3A",
    315 => X"3B",
    316 => X"3C",
    317 => X"3D",
    318 => X"3E",
    319 => X"3F",
    320 => X"40",
    321 => X"41",
    322 => X"42",
    323 => X"43",
    324 => X"44",
    325 => X"45",
    326 => X"46",
    327 => X"47",
    328 => X"48",
    329 => X"49",
    330 => X"4A",
    331 => X"4B",
    332 => X"4C",
    333 => X"4D",
    334 => X"4E",
    335 => X"4F",
    336 => X"50",
    337 => X"51",
    338 => X"52",
    339 => X"53",
    340 => X"54",
    341 => X"55",
    342 => X"56",
    343 => X"57",
    344 => X"58",
    345 => X"59",
    346 => X"5A",
    347 => X"5B",
    348 => X"5C",
    349 => X"5D",
    350 => X"5E",
    351 => X"5F",
    352 => X"60",
    353 => X"61",
    354 => X"62",
    355 => X"63",
    356 => X"64",
    357 => X"65",
    358 => X"66",
    359 => X"67",
    360 => X"68",
    361 => X"69",
    362 => X"6A",
    363 => X"6B",
    364 => X"6C",
    365 => X"6D",
    366 => X"6E",
    367 => X"6F",
    368 => X"70",
    369 => X"71",
    370 => X"72",
    371 => X"73",
    372 => X"74",
    373 => X"75",
    374 => X"76",
    375 => X"77",
    376 => X"78",
    377 => X"79",
    378 => X"7A",
    379 => X"7B",
    380 => X"7C",
    381 => X"7D",
    382 => X"7E",
    383 => X"7F",
    384 => X"80",
    385 => X"81",
    386 => X"82",
    387 => X"83",
    388 => X"84",
    389 => X"85",
    390 => X"86",
    391 => X"87",
    392 => X"88",
    393 => X"89",
    394 => X"8A",
    395 => X"8B",
    396 => X"8C",
    397 => X"8D",
    398 => X"8E",
    399 => X"8F",
    400 => X"90",
    401 => X"91",
    402 => X"92",
    403 => X"93",
    404 => X"94",
    405 => X"95",
    406 => X"96",
    407 => X"97",
    408 => X"98",
    409 => X"99",
    410 => X"9A",
    411 => X"9B",
    412 => X"9C",
    413 => X"9D",
    414 => X"9E",
    415 => X"9F",
    416 => X"A0",
    417 => X"A1",
    418 => X"A2",
    419 => X"A3",
    420 => X"A4",
    421 => X"A5",
    422 => X"A6",
    423 => X"A7",
    424 => X"A8",
    425 => X"A9",
    426 => X"AA",
    427 => X"AB",
    428 => X"AC",
    429 => X"AD",
    430 => X"AE",
    431 => X"AF",
    432 => X"B0",
    433 => X"B1",
    434 => X"B2",
    435 => X"B3",
    436 => X"B4",
    437 => X"B5",
    438 => X"B6",
    439 => X"B7",
    440 => X"B8",
    441 => X"B9",
    442 => X"BA",
    443 => X"BB",
    444 => X"BC",
    445 => X"BD",
    446 => X"BE",
    447 => X"BF",
    448 => X"C0",
    449 => X"C1",
    450 => X"C2",
    451 => X"C3",
    452 => X"C4",
    453 => X"C5",
    454 => X"C6",
    455 => X"C7",
    456 => X"C8",
    457 => X"C9",
    458 => X"CA",
    459 => X"CB",
    460 => X"CC",
    461 => X"CD",
    462 => X"CE",
    463 => X"CF",
    464 => X"D0",
    465 => X"D1",
    466 => X"D2",
    467 => X"D3",
    468 => X"D4",
    469 => X"D5",
    470 => X"D6",
    471 => X"D7",
    472 => X"D8",
    473 => X"D9",
    474 => X"DA",
    475 => X"DB",
    476 => X"DC",
    477 => X"DD",
    478 => X"DE",
    479 => X"DF",
    480 => X"E0",
    481 => X"E1",
    482 => X"E2",
    483 => X"E3",
    484 => X"E4",
    485 => X"E5",
    486 => X"E6",
    487 => X"E7",
    488 => X"E8",
    489 => X"E9",
    490 => X"EA",
    491 => X"EB",
    492 => X"EC",
    493 => X"ED",
    494 => X"EE",
    495 => X"EF",
    496 => X"F0",
    497 => X"F1",
    498 => X"F2",
    499 => X"F3",
    500 => X"F4",
    501 => X"F5",
    502 => X"F6",
    503 => X"F7",
    504 => X"F8",
    505 => X"F9",
    506 => X"FA",
    507 => X"FB",
    508 => X"FC",
    509 => X"FD",
    510 => X"FE",
    511 => X"FF",
    512 => X"00",
    513 => X"01",
    514 => X"02",
    515 => X"03",
    516 => X"04",
    517 => X"05",
    518 => X"06",
    519 => X"07",
    520 => X"08",
    521 => X"09",
    522 => X"0A",
    523 => X"0B",
    524 => X"0C",
    525 => X"0D",
    526 => X"0E",
    527 => X"0F",
    528 => X"10",
    529 => X"11",
    530 => X"12",
    531 => X"13",
    532 => X"14",
    533 => X"15",
    534 => X"16",
    535 => X"17",
    536 => X"18",
    537 => X"19",
    538 => X"1A",
    539 => X"1B",
    540 => X"1C",
    541 => X"1D",
    542 => X"1E",
    543 => X"1F",
    544 => X"20",
    545 => X"21",
    546 => X"22",
    547 => X"23",
    548 => X"24",
    549 => X"25",
    550 => X"26",
    551 => X"27",
    552 => X"28",
    553 => X"29",
    554 => X"2A",
    555 => X"2B",
    556 => X"2C",
    557 => X"2D",
    558 => X"2E",
    559 => X"2F",
    560 => X"30",
    561 => X"31",
    562 => X"32",
    563 => X"33",
    564 => X"34",
    565 => X"35",
    566 => X"36",
    567 => X"37",
    568 => X"38",
    569 => X"39",
    570 => X"3A",
    571 => X"3B",
    572 => X"3C",
    573 => X"3D",
    574 => X"3E",
    575 => X"3F",
    576 => X"40",
    577 => X"41",
    578 => X"42",
    579 => X"43",
    580 => X"44",
    581 => X"45",
    582 => X"46",
    583 => X"47",
    584 => X"48",
    585 => X"49",
    586 => X"4A",
    587 => X"4B",
    588 => X"4C",
    589 => X"4D",
    590 => X"4E",
    591 => X"4F",
    592 => X"50",
    593 => X"51",
    594 => X"52",
    595 => X"53",
    596 => X"54",
    597 => X"55",
    598 => X"56",
    599 => X"57",
    600 => X"58",
    601 => X"59",
    602 => X"5A",
    603 => X"5B",
    604 => X"5C",
    605 => X"5D",
    606 => X"5E",
    607 => X"5F",
    608 => X"60",
    609 => X"61",
    610 => X"62",
    611 => X"63",
    612 => X"64",
    613 => X"65",
    614 => X"66",
    615 => X"67",
    616 => X"68",
    617 => X"69",
    618 => X"6A",
    619 => X"6B",
    620 => X"6C",
    621 => X"6D",
    622 => X"6E",
    623 => X"6F",
    624 => X"70",
    625 => X"71",
    626 => X"72",
    627 => X"73",
    628 => X"74",
    629 => X"75",
    630 => X"76",
    631 => X"77",
    632 => X"78",
    633 => X"79",
    634 => X"7A",
    635 => X"7B",
    636 => X"7C",
    637 => X"7D",
    638 => X"7E",
    639 => X"7F",
    640 => X"80",
    641 => X"81",
    642 => X"82",
    643 => X"83",
    644 => X"84",
    645 => X"85",
    646 => X"86",
    647 => X"87",
    648 => X"88",
    649 => X"89",
    650 => X"8A",
    651 => X"8B",
    652 => X"8C",
    653 => X"8D",
    654 => X"8E",
    655 => X"8F",
    656 => X"90",
    657 => X"91",
    658 => X"92",
    659 => X"93",
    660 => X"94",
    661 => X"95",
    662 => X"96",
    663 => X"97",
    664 => X"98",
    665 => X"99",
    666 => X"9A",
    667 => X"9B",
    668 => X"9C",
    669 => X"9D",
    670 => X"9E",
    671 => X"9F",
    672 => X"A0",
    673 => X"A1",
    674 => X"A2",
    675 => X"A3",
    676 => X"A4",
    677 => X"A5",
    678 => X"A6",
    679 => X"A7",
    680 => X"A8",
    681 => X"A9",
    682 => X"AA",
    683 => X"AB",
    684 => X"AC",
    685 => X"AD",
    686 => X"AE",
    687 => X"AF",
    688 => X"B0",
    689 => X"B1",
    690 => X"B2",
    691 => X"B3",
    692 => X"B4",
    693 => X"B5",
    694 => X"B6",
    695 => X"B7",
    696 => X"B8",
    697 => X"B9",
    698 => X"BA",
    699 => X"BB",
    700 => X"BC",
    701 => X"BD",
    702 => X"BE",
    703 => X"BF",
    704 => X"C0",
    705 => X"C1",
    706 => X"C2",
    707 => X"C3",
    708 => X"C4",
    709 => X"C5",
    710 => X"C6",
    711 => X"C7",
    712 => X"C8",
    713 => X"C9",
    714 => X"CA",
    715 => X"CB",
    716 => X"CC",
    717 => X"CD",
    718 => X"CE",
    719 => X"CF",
    720 => X"D0",
    721 => X"D1",
    722 => X"D2",
    723 => X"D3",
    724 => X"D4",
    725 => X"D5",
    726 => X"D6",
    727 => X"D7",
    728 => X"D8",
    729 => X"D9",
    730 => X"DA",
    731 => X"DB",
    732 => X"DC",
    733 => X"DD",
    734 => X"DE",
    735 => X"DF",
    736 => X"E0",
    737 => X"E1",
    738 => X"E2",
    739 => X"E3",
    740 => X"E4",
    741 => X"E5",
    742 => X"E6",
    743 => X"E7",
    744 => X"E8",
    745 => X"E9",
    746 => X"EA",
    747 => X"EB",
    748 => X"EC",
    749 => X"ED",
    750 => X"EE",
    751 => X"EF",
    752 => X"F0",
    753 => X"F1",
    754 => X"F2",
    755 => X"F3",
    756 => X"F4",
    757 => X"F5",
    758 => X"F6",
    759 => X"F7",
    760 => X"F8",
    761 => X"F9",
    762 => X"FA",
    763 => X"FB",
    764 => X"FC",
    765 => X"FD",
    766 => X"FE",
    767 => X"FF",
    768 => X"00",
    769 => X"01",
    770 => X"02",
    771 => X"03",
    772 => X"04",
    773 => X"05",
    774 => X"06",
    775 => X"07",
    776 => X"08",
    777 => X"09",
    778 => X"0A",
    779 => X"0B",
    780 => X"0C",
    781 => X"0D",
    782 => X"0E",
    783 => X"0F",
    784 => X"10",
    785 => X"11",
    786 => X"12",
    787 => X"13",
    788 => X"14",
    789 => X"15",
    790 => X"16",
    791 => X"17",
    792 => X"18",
    793 => X"19",
    794 => X"1A",
    795 => X"1B",
    796 => X"1C",
    797 => X"1D",
    798 => X"1E",
    799 => X"1F",
    800 => X"20",
    801 => X"21",
    802 => X"22",
    803 => X"23",
    804 => X"24",
    805 => X"25",
    806 => X"26",
    807 => X"27",
    808 => X"28",
    809 => X"29",
    810 => X"2A",
    811 => X"2B",
    812 => X"2C",
    813 => X"2D",
    814 => X"2E",
    815 => X"2F",
    816 => X"30",
    817 => X"31",
    818 => X"32",
    819 => X"33",
    820 => X"34",
    821 => X"35",
    822 => X"36",
    823 => X"37",
    824 => X"38",
    825 => X"39",
    826 => X"3A",
    827 => X"3B",
    828 => X"3C",
    829 => X"3D",
    830 => X"3E",
    831 => X"3F",
    832 => X"40",
    833 => X"41",
    834 => X"42",
    835 => X"43",
    836 => X"44",
    837 => X"45",
    838 => X"46",
    839 => X"47",
    840 => X"48",
    841 => X"49",
    842 => X"4A",
    843 => X"4B",
    844 => X"4C",
    845 => X"4D",
    846 => X"4E",
    847 => X"4F",
    848 => X"50",
    849 => X"51",
    850 => X"52",
    851 => X"53",
    852 => X"54",
    853 => X"55",
    854 => X"56",
    855 => X"57",
    856 => X"58",
    857 => X"59",
    858 => X"5A",
    859 => X"5B",
    860 => X"5C",
    861 => X"5D",
    862 => X"5E",
    863 => X"5F",
    864 => X"60",
    865 => X"61",
    866 => X"62",
    867 => X"63",
    868 => X"64",
    869 => X"65",
    870 => X"66",
    871 => X"67",
    872 => X"68",
    873 => X"69",
    874 => X"6A",
    875 => X"6B",
    876 => X"6C",
    877 => X"6D",
    878 => X"6E",
    879 => X"6F",
    880 => X"70",
    881 => X"71",
    882 => X"72",
    883 => X"73",
    884 => X"74",
    885 => X"75",
    886 => X"76",
    887 => X"77",
    888 => X"78",
    889 => X"79",
    890 => X"7A",
    891 => X"7B",
    892 => X"7C",
    893 => X"7D",
    894 => X"7E",
    895 => X"7F",
    896 => X"80",
    897 => X"81",
    898 => X"82",
    899 => X"83",
    900 => X"84",
    901 => X"85",
    902 => X"86",
    903 => X"87",
    904 => X"88",
    905 => X"89",
    906 => X"8A",
    907 => X"8B",
    908 => X"8C",
    909 => X"8D",
    910 => X"8E",
    911 => X"8F",
    912 => X"90",
    913 => X"91",
    914 => X"92",
    915 => X"93",
    916 => X"94",
    917 => X"95",
    918 => X"96",
    919 => X"97",
    920 => X"98",
    921 => X"99",
    922 => X"9A",
    923 => X"9B",
    924 => X"9C",
    925 => X"9D",
    926 => X"9E",
    927 => X"9F",
    928 => X"A0",
    929 => X"A1",
    930 => X"A2",
    931 => X"A3",
    932 => X"A4",
    933 => X"A5",
    934 => X"A6",
    935 => X"A7",
    936 => X"A8",
    937 => X"A9",
    938 => X"AA",
    939 => X"AB",
    940 => X"AC",
    941 => X"AD",
    942 => X"AE",
    943 => X"AF",
    944 => X"B0",
    945 => X"B1",
    946 => X"B2",
    947 => X"B3",
    948 => X"B4",
    949 => X"B5",
    950 => X"B6",
    951 => X"B7",
    952 => X"B8",
    953 => X"B9",
    954 => X"BA",
    955 => X"BB",
    956 => X"BC",
    957 => X"BD",
    958 => X"BE",
    959 => X"BF",
    960 => X"C0",
    961 => X"C1",
    962 => X"C2",
    963 => X"C3",
    964 => X"C4",
    965 => X"C5",
    966 => X"C6",
    967 => X"C7",
    968 => X"C8",
    969 => X"C9",
    970 => X"CA",
    971 => X"CB",
    972 => X"CC",
    973 => X"CD",
    974 => X"CE",
    975 => X"CF",
    976 => X"D0",
    977 => X"D1",
    978 => X"D2",
    979 => X"D3",
    980 => X"D4",
    981 => X"D5",
    982 => X"D6",
    983 => X"D7",
    984 => X"D8",
    985 => X"D9",
    986 => X"DA",
    987 => X"DB",
    988 => X"DC",
    989 => X"DD",
    990 => X"DE",
    991 => X"DF",
    992 => X"E0",
    993 => X"E1",
    994 => X"E2",
    995 => X"E3",
    996 => X"E4",
    997 => X"E5",
    998 => X"E6",
    999 => X"E7",
    1000 => X"E8",
    1001 => X"E9",
    1002 => X"EA",
    1003 => X"EB",
    1004 => X"EC",
    1005 => X"ED",
    1006 => X"EE",
    1007 => X"EF",
    1008 => X"F0",
    1009 => X"F1",
    1010 => X"F2",
    1011 => X"F3",
    1012 => X"F4",
    1013 => X"F5",
    1014 => X"F6",
    1015 => X"F7",
    1016 => X"F8",
    1017 => X"F9",
    1018 => X"FA",
    1019 => X"FB",
    1020 => X"FC",
    1021 => X"FD",
    1022 => X"FE",
    1023 => X"FF",
    1024 => X"00",
    1025 => X"01",
    1026 => X"02",
    1027 => X"03",
    1028 => X"04",
    1029 => X"05",
    1030 => X"06",
    1031 => X"07",
    1032 => X"08",
    1033 => X"09",
    1034 => X"0A",
    1035 => X"0B",
    1036 => X"0C",
    1037 => X"0D",
    1038 => X"0E",
    1039 => X"0F",
    1040 => X"10",
    1041 => X"11",
    1042 => X"12",
    1043 => X"13",
    1044 => X"14",
    1045 => X"15",
    1046 => X"16",
    1047 => X"17",
    1048 => X"18",
    1049 => X"19",
    1050 => X"1A",
    1051 => X"1B",
    1052 => X"1C",
    1053 => X"1D",
    1054 => X"1E",
    1055 => X"1F",
    1056 => X"20",
    1057 => X"21",
    1058 => X"22",
    1059 => X"23",
    1060 => X"24",
    1061 => X"25",
    1062 => X"26",
    1063 => X"27",
    1064 => X"28",
    1065 => X"29",
    1066 => X"2A",
    1067 => X"2B",
    1068 => X"2C",
    1069 => X"2D",
    1070 => X"2E",
    1071 => X"2F",
    1072 => X"30",
    1073 => X"31",
    1074 => X"32",
    1075 => X"33",
    1076 => X"34",
    1077 => X"35",
    1078 => X"36",
    1079 => X"37",
    1080 => X"38",
    1081 => X"39",
    1082 => X"3A",
    1083 => X"3B",
    1084 => X"3C",
    1085 => X"3D",
    1086 => X"3E",
    1087 => X"3F",
    1088 => X"40",
    1089 => X"41",
    1090 => X"42",
    1091 => X"43",
    1092 => X"44",
    1093 => X"45",
    1094 => X"46",
    1095 => X"47",
    1096 => X"48",
    1097 => X"49",
    1098 => X"4A",
    1099 => X"4B",
    1100 => X"4C",
    1101 => X"4D",
    1102 => X"4E",
    1103 => X"4F",
    1104 => X"50",
    1105 => X"51",
    1106 => X"52",
    1107 => X"53",
    1108 => X"54",
    1109 => X"55",
    1110 => X"56",
    1111 => X"57",
    1112 => X"58",
    1113 => X"59",
    1114 => X"5A",
    1115 => X"5B",
    1116 => X"5C",
    1117 => X"5D",
    1118 => X"5E",
    1119 => X"5F",
    1120 => X"60",
    1121 => X"61",
    1122 => X"62",
    1123 => X"63",
    1124 => X"64",
    1125 => X"65",
    1126 => X"66",
    1127 => X"67",
    1128 => X"68",
    1129 => X"69",
    1130 => X"6A",
    1131 => X"6B",
    1132 => X"6C",
    1133 => X"6D",
    1134 => X"6E",
    1135 => X"6F",
    1136 => X"70",
    1137 => X"71",
    1138 => X"72",
    1139 => X"73",
    1140 => X"74",
    1141 => X"75",
    1142 => X"76",
    1143 => X"77",
    1144 => X"78",
    1145 => X"79",
    1146 => X"7A",
    1147 => X"7B",
    1148 => X"7C",
    1149 => X"7D",
    1150 => X"7E",
    1151 => X"7F",
    1152 => X"80",
    1153 => X"81",
    1154 => X"82",
    1155 => X"83",
    1156 => X"84",
    1157 => X"85",
    1158 => X"86",
    1159 => X"87",
    1160 => X"88",
    1161 => X"89",
    1162 => X"8A",
    1163 => X"8B",
    1164 => X"8C",
    1165 => X"8D",
    1166 => X"8E",
    1167 => X"8F",
    1168 => X"90",
    1169 => X"91",
    1170 => X"92",
    1171 => X"93",
    1172 => X"94",
    1173 => X"95",
    1174 => X"96",
    1175 => X"97",
    1176 => X"98",
    1177 => X"99",
    1178 => X"9A",
    1179 => X"9B",
    1180 => X"9C",
    1181 => X"9D",
    1182 => X"9E",
    1183 => X"9F",
    1184 => X"A0",
    1185 => X"A1",
    1186 => X"A2",
    1187 => X"A3",
    1188 => X"A4",
    1189 => X"A5",
    1190 => X"A6",
    1191 => X"A7",
    1192 => X"A8",
    1193 => X"A9",
    1194 => X"AA",
    1195 => X"AB",
    1196 => X"AC",
    1197 => X"AD",
    1198 => X"AE",
    1199 => X"AF",
    1200 => X"B0",
    1201 => X"B1",
    1202 => X"B2",
    1203 => X"B3",
    1204 => X"B4",
    1205 => X"B5",
    1206 => X"B6",
    1207 => X"B7",
    1208 => X"B8",
    1209 => X"B9",
    1210 => X"BA",
    1211 => X"BB",
    1212 => X"BC",
    1213 => X"BD",
    1214 => X"BE",
    1215 => X"BF",
    1216 => X"C0",
    1217 => X"C1",
    1218 => X"C2",
    1219 => X"C3",
    1220 => X"C4",
    1221 => X"C5",
    1222 => X"C6",
    1223 => X"C7",
    1224 => X"C8",
    1225 => X"C9",
    1226 => X"CA",
    1227 => X"CB",
    1228 => X"CC",
    1229 => X"CD",
    1230 => X"CE",
    1231 => X"CF",
    1232 => X"D0",
    1233 => X"D1",
    1234 => X"D2",
    1235 => X"D3",
    1236 => X"D4",
    1237 => X"D5",
    1238 => X"D6",
    1239 => X"D7",
    1240 => X"D8",
    1241 => X"D9",
    1242 => X"DA",
    1243 => X"DB",
    1244 => X"DC",
    1245 => X"DD",
    1246 => X"DE",
    1247 => X"DF",
    1248 => X"E0",
    1249 => X"E1",
    1250 => X"E2",
    1251 => X"E3",
    1252 => X"E4",
    1253 => X"E5",
    1254 => X"E6",
    1255 => X"E7",
    1256 => X"E8",
    1257 => X"E9",
    1258 => X"EA",
    1259 => X"EB",
    1260 => X"EC",
    1261 => X"ED",
    1262 => X"EE",
    1263 => X"EF",
    1264 => X"F0",
    1265 => X"F1",
    1266 => X"F2",
    1267 => X"F3",
    1268 => X"F4",
    1269 => X"F5",
    1270 => X"F6",
    1271 => X"F7",
    1272 => X"F8",
    1273 => X"F9",
    1274 => X"FA",
    1275 => X"FB",
    1276 => X"FC",
    1277 => X"FD",
    1278 => X"FE",
    1279 => X"FF",
    1280 => X"00",
    1281 => X"01",
    1282 => X"02",
    1283 => X"03",
    1284 => X"04",
    1285 => X"05",
    1286 => X"06",
    1287 => X"07",
    1288 => X"08",
    1289 => X"09",
    1290 => X"0A",
    1291 => X"0B",
    1292 => X"0C",
    1293 => X"0D",
    1294 => X"0E",
    1295 => X"0F",
    1296 => X"10",
    1297 => X"11",
    1298 => X"12",
    1299 => X"13",
    1300 => X"14",
    1301 => X"15",
    1302 => X"16",
    1303 => X"17",
    1304 => X"18",
    1305 => X"19",
    1306 => X"1A",
    1307 => X"1B",
    1308 => X"1C",
    1309 => X"1D",
    1310 => X"1E",
    1311 => X"1F",
    1312 => X"20",
    1313 => X"21",
    1314 => X"22",
    1315 => X"23",
    1316 => X"24",
    1317 => X"25",
    1318 => X"26",
    1319 => X"27",
    1320 => X"28",
    1321 => X"29",
    1322 => X"2A",
    1323 => X"2B",
    1324 => X"2C",
    1325 => X"2D",
    1326 => X"2E",
    1327 => X"2F",
    1328 => X"30",
    1329 => X"31",
    1330 => X"32",
    1331 => X"33",
    1332 => X"34",
    1333 => X"35",
    1334 => X"36",
    1335 => X"37",
    1336 => X"38",
    1337 => X"39",
    1338 => X"3A",
    1339 => X"3B",
    1340 => X"3C",
    1341 => X"3D",
    1342 => X"3E",
    1343 => X"3F",
    1344 => X"40",
    1345 => X"41",
    1346 => X"42",
    1347 => X"43",
    1348 => X"44",
    1349 => X"45",
    1350 => X"46",
    1351 => X"47",
    1352 => X"48",
    1353 => X"49",
    1354 => X"4A",
    1355 => X"4B",
    1356 => X"4C",
    1357 => X"4D",
    1358 => X"4E",
    1359 => X"4F",
    1360 => X"50",
    1361 => X"51",
    1362 => X"52",
    1363 => X"53",
    1364 => X"54",
    1365 => X"55",
    1366 => X"56",
    1367 => X"57",
    1368 => X"58",
    1369 => X"59",
    1370 => X"5A",
    1371 => X"5B",
    1372 => X"5C",
    1373 => X"5D",
    1374 => X"5E",
    1375 => X"5F",
    1376 => X"60",
    1377 => X"61",
    1378 => X"62",
    1379 => X"63",
    1380 => X"64",
    1381 => X"65",
    1382 => X"66",
    1383 => X"67",
    1384 => X"68",
    1385 => X"69",
    1386 => X"6A",
    1387 => X"6B",
    1388 => X"6C",
    1389 => X"6D",
    1390 => X"6E",
    1391 => X"6F",
    1392 => X"70",
    1393 => X"71",
    1394 => X"72",
    1395 => X"73",
    1396 => X"74",
    1397 => X"75",
    1398 => X"76",
    1399 => X"77",
    1400 => X"78",
    1401 => X"79",
    1402 => X"7A",
    1403 => X"7B",
    1404 => X"7C",
    1405 => X"7D",
    1406 => X"7E",
    1407 => X"7F",
    1408 => X"80",
    1409 => X"81",
    1410 => X"82",
    1411 => X"83",
    1412 => X"84",
    1413 => X"85",
    1414 => X"86",
    1415 => X"87",
    1416 => X"88",
    1417 => X"89",
    1418 => X"8A",
    1419 => X"8B",
    1420 => X"8C",
    1421 => X"8D",
    1422 => X"8E",
    1423 => X"8F",
    1424 => X"90",
    1425 => X"91",
    1426 => X"92",
    1427 => X"93",
    1428 => X"94",
    1429 => X"95",
    1430 => X"96",
    1431 => X"97",
    1432 => X"98",
    1433 => X"99",
    1434 => X"9A",
    1435 => X"9B",
    1436 => X"9C",
    1437 => X"9D",
    1438 => X"9E",
    1439 => X"9F",
    1440 => X"A0",
    1441 => X"A1",
    1442 => X"A2",
    1443 => X"A3",
    1444 => X"A4",
    1445 => X"A5",
    1446 => X"A6",
    1447 => X"A7",
    1448 => X"A8",
    1449 => X"A9",
    1450 => X"AA",
    1451 => X"AB",
    1452 => X"AC",
    1453 => X"AD",
    1454 => X"AE",
    1455 => X"AF",
    1456 => X"B0",
    1457 => X"B1",
    1458 => X"B2",
    1459 => X"B3",
    1460 => X"B4",
    1461 => X"B5",
    1462 => X"B6",
    1463 => X"B7",
    1464 => X"B8",
    1465 => X"B9",
    1466 => X"BA",
    1467 => X"BB",
    1468 => X"BC",
    1469 => X"BD",
    1470 => X"BE",
    1471 => X"BF",
    1472 => X"C0",
    1473 => X"C1",
    1474 => X"C2",
    1475 => X"C3",
    1476 => X"C4",
    1477 => X"C5",
    1478 => X"C6",
    1479 => X"C7",
    1480 => X"C8",
    1481 => X"C9",
    1482 => X"CA",
    1483 => X"CB",
    1484 => X"CC",
    1485 => X"CD",
    1486 => X"CE",
    1487 => X"CF",
    1488 => X"D0",
    1489 => X"D1",
    1490 => X"D2",
    1491 => X"D3",
    1492 => X"D4",
    1493 => X"D5",
    1494 => X"D6",
    1495 => X"D7",
    1496 => X"D8",
    1497 => X"D9",
    1498 => X"DA",
    1499 => X"DB",
    1500 => X"DC",
    1501 => X"DD",
    1502 => X"DE",
    1503 => X"DF",
    1504 => X"E0",
    1505 => X"E1",
    1506 => X"E2",
    1507 => X"E3",
    1508 => X"E4",
    1509 => X"E5",
    1510 => X"E6",
    1511 => X"E7",
    1512 => X"E8",
    1513 => X"E9",
    1514 => X"EA",
    1515 => X"EB",
    1516 => X"EC",
    1517 => X"ED",
    1518 => X"EE",
    1519 => X"EF",
    1520 => X"F0",
    1521 => X"F1",
    1522 => X"F2",
    1523 => X"F3",
    1524 => X"F4",
    1525 => X"F5",
    1526 => X"F6",
    1527 => X"F7",
    1528 => X"F8",
    1529 => X"F9",
    1530 => X"FA",
    1531 => X"FB",
    1532 => X"FC",
    1533 => X"FD",
    1534 => X"FE",
    1535 => X"FF",
    1536 => X"00",
    1537 => X"01",
    1538 => X"02",
    1539 => X"03",
    1540 => X"04",
    1541 => X"05",
    1542 => X"06",
    1543 => X"07",
    1544 => X"08",
    1545 => X"09",
    1546 => X"0A",
    1547 => X"0B",
    1548 => X"0C",
    1549 => X"0D",
    1550 => X"0E",
    1551 => X"0F",
    1552 => X"10",
    1553 => X"11",
    1554 => X"12",
    1555 => X"13",
    1556 => X"14",
    1557 => X"15",
    1558 => X"16",
    1559 => X"17",
    1560 => X"18",
    1561 => X"19",
    1562 => X"1A",
    1563 => X"1B",
    1564 => X"1C",
    1565 => X"1D",
    1566 => X"1E",
    1567 => X"1F",
    1568 => X"20",
    1569 => X"21",
    1570 => X"22",
    1571 => X"23",
    1572 => X"24",
    1573 => X"25",
    1574 => X"26",
    1575 => X"27",
    1576 => X"28",
    1577 => X"29",
    1578 => X"2A",
    1579 => X"2B",
    1580 => X"2C",
    1581 => X"2D",
    1582 => X"2E",
    1583 => X"2F",
    1584 => X"30",
    1585 => X"31",
    1586 => X"32",
    1587 => X"33",
    1588 => X"34",
    1589 => X"35",
    1590 => X"36",
    1591 => X"37",
    1592 => X"38",
    1593 => X"39",
    1594 => X"3A",
    1595 => X"3B",
    1596 => X"3C",
    1597 => X"3D",
    1598 => X"3E",
    1599 => X"3F",
    1600 => X"40",
    1601 => X"41",
    1602 => X"42",
    1603 => X"43",
    1604 => X"44",
    1605 => X"45",
    1606 => X"46",
    1607 => X"47",
    1608 => X"48",
    1609 => X"49",
    1610 => X"4A",
    1611 => X"4B",
    1612 => X"4C",
    1613 => X"4D",
    1614 => X"4E",
    1615 => X"4F",
    1616 => X"50",
    1617 => X"51",
    1618 => X"52",
    1619 => X"53",
    1620 => X"54",
    1621 => X"55",
    1622 => X"56",
    1623 => X"57",
    1624 => X"58",
    1625 => X"59",
    1626 => X"5A",
    1627 => X"5B",
    1628 => X"5C",
    1629 => X"5D",
    1630 => X"5E",
    1631 => X"5F",
    1632 => X"60",
    1633 => X"61",
    1634 => X"62",
    1635 => X"63",
    1636 => X"64",
    1637 => X"65",
    1638 => X"66",
    1639 => X"67",
    1640 => X"68",
    1641 => X"69",
    1642 => X"6A",
    1643 => X"6B",
    1644 => X"6C",
    1645 => X"6D",
    1646 => X"6E",
    1647 => X"6F",
    1648 => X"70",
    1649 => X"71",
    1650 => X"72",
    1651 => X"73",
    1652 => X"74",
    1653 => X"75",
    1654 => X"76",
    1655 => X"77",
    1656 => X"78",
    1657 => X"79",
    1658 => X"7A",
    1659 => X"7B",
    1660 => X"7C",
    1661 => X"7D",
    1662 => X"7E",
    1663 => X"7F",
    1664 => X"80",
    1665 => X"81",
    1666 => X"82",
    1667 => X"83",
    1668 => X"84",
    1669 => X"85",
    1670 => X"86",
    1671 => X"87",
    1672 => X"88",
    1673 => X"89",
    1674 => X"8A",
    1675 => X"8B",
    1676 => X"8C",
    1677 => X"8D",
    1678 => X"8E",
    1679 => X"8F",
    1680 => X"90",
    1681 => X"91",
    1682 => X"92",
    1683 => X"93",
    1684 => X"94",
    1685 => X"95",
    1686 => X"96",
    1687 => X"97",
    1688 => X"98",
    1689 => X"99",
    1690 => X"9A",
    1691 => X"9B",
    1692 => X"9C",
    1693 => X"9D",
    1694 => X"9E",
    1695 => X"9F",
    1696 => X"A0",
    1697 => X"A1",
    1698 => X"A2",
    1699 => X"A3",
    1700 => X"A4",
    1701 => X"A5",
    1702 => X"A6",
    1703 => X"A7",
    1704 => X"A8",
    1705 => X"A9",
    1706 => X"AA",
    1707 => X"AB",
    1708 => X"AC",
    1709 => X"AD",
    1710 => X"AE",
    1711 => X"AF",
    1712 => X"B0",
    1713 => X"B1",
    1714 => X"B2",
    1715 => X"B3",
    1716 => X"B4",
    1717 => X"B5",
    1718 => X"B6",
    1719 => X"B7",
    1720 => X"B8",
    1721 => X"B9",
    1722 => X"BA",
    1723 => X"BB",
    1724 => X"BC",
    1725 => X"BD",
    1726 => X"BE",
    1727 => X"BF",
    1728 => X"C0",
    1729 => X"C1",
    1730 => X"C2",
    1731 => X"C3",
    1732 => X"C4",
    1733 => X"C5",
    1734 => X"C6",
    1735 => X"C7",
    1736 => X"C8",
    1737 => X"C9",
    1738 => X"CA",
    1739 => X"CB",
    1740 => X"CC",
    1741 => X"CD",
    1742 => X"CE",
    1743 => X"CF",
    1744 => X"D0",
    1745 => X"D1",
    1746 => X"D2",
    1747 => X"D3",
    1748 => X"D4",
    1749 => X"D5",
    1750 => X"D6",
    1751 => X"D7",
    1752 => X"D8",
    1753 => X"D9",
    1754 => X"DA",
    1755 => X"DB",
    1756 => X"DC",
    1757 => X"DD",
    1758 => X"DE",
    1759 => X"DF",
    1760 => X"E0",
    1761 => X"E1",
    1762 => X"E2",
    1763 => X"E3",
    1764 => X"E4",
    1765 => X"E5",
    1766 => X"E6",
    1767 => X"E7",
    1768 => X"E8",
    1769 => X"E9",
    1770 => X"EA",
    1771 => X"EB",
    1772 => X"EC",
    1773 => X"ED",
    1774 => X"EE",
    1775 => X"EF",
    1776 => X"F0",
    1777 => X"F1",
    1778 => X"F2",
    1779 => X"F3",
    1780 => X"F4",
    1781 => X"F5",
    1782 => X"F6",
    1783 => X"F7",
    1784 => X"F8",
    1785 => X"F9",
    1786 => X"FA",
    1787 => X"FB",
    1788 => X"FC",
    1789 => X"FD",
    1790 => X"FE",
    1791 => X"FF",
    1792 => X"00",
    1793 => X"01",
    1794 => X"02",
    1795 => X"03",
    1796 => X"04",
    1797 => X"05",
    1798 => X"06",
    1799 => X"07",
    1800 => X"08",
    1801 => X"09",
    1802 => X"0A",
    1803 => X"0B",
    1804 => X"0C",
    1805 => X"0D",
    1806 => X"0E",
    1807 => X"0F",
    1808 => X"10",
    1809 => X"11",
    1810 => X"12",
    1811 => X"13",
    1812 => X"14",
    1813 => X"15",
    1814 => X"16",
    1815 => X"17",
    1816 => X"18",
    1817 => X"19",
    1818 => X"1A",
    1819 => X"1B",
    1820 => X"1C",
    1821 => X"1D",
    1822 => X"1E",
    1823 => X"1F",
    1824 => X"20",
    1825 => X"21",
    1826 => X"22",
    1827 => X"23",
    1828 => X"24",
    1829 => X"25",
    1830 => X"26",
    1831 => X"27",
    1832 => X"28",
    1833 => X"29",
    1834 => X"2A",
    1835 => X"2B",
    1836 => X"2C",
    1837 => X"2D",
    1838 => X"2E",
    1839 => X"2F",
    1840 => X"30",
    1841 => X"31",
    1842 => X"32",
    1843 => X"33",
    1844 => X"34",
    1845 => X"35",
    1846 => X"36",
    1847 => X"37",
    1848 => X"38",
    1849 => X"39",
    1850 => X"3A",
    1851 => X"3B",
    1852 => X"3C",
    1853 => X"3D",
    1854 => X"3E",
    1855 => X"3F",
    1856 => X"40",
    1857 => X"41",
    1858 => X"42",
    1859 => X"43",
    1860 => X"44",
    1861 => X"45",
    1862 => X"46",
    1863 => X"47",
    1864 => X"48",
    1865 => X"49",
    1866 => X"4A",
    1867 => X"4B",
    1868 => X"4C",
    1869 => X"4D",
    1870 => X"4E",
    1871 => X"4F",
    1872 => X"50",
    1873 => X"51",
    1874 => X"52",
    1875 => X"53",
    1876 => X"54",
    1877 => X"55",
    1878 => X"56",
    1879 => X"57",
    1880 => X"58",
    1881 => X"59",
    1882 => X"5A",
    1883 => X"5B",
    1884 => X"5C",
    1885 => X"5D",
    1886 => X"5E",
    1887 => X"5F",
    1888 => X"60",
    1889 => X"61",
    1890 => X"62",
    1891 => X"63",
    1892 => X"64",
    1893 => X"65",
    1894 => X"66",
    1895 => X"67",
    1896 => X"68",
    1897 => X"69",
    1898 => X"6A",
    1899 => X"6B",
    1900 => X"6C",
    1901 => X"6D",
    1902 => X"6E",
    1903 => X"6F",
    1904 => X"70",
    1905 => X"71",
    1906 => X"72",
    1907 => X"73",
    1908 => X"74",
    1909 => X"75",
    1910 => X"76",
    1911 => X"77",
    1912 => X"78",
    1913 => X"79",
    1914 => X"7A",
    1915 => X"7B",
    1916 => X"7C",
    1917 => X"7D",
    1918 => X"7E",
    1919 => X"7F",
    1920 => X"80",
    1921 => X"81",
    1922 => X"82",
    1923 => X"83",
    1924 => X"84",
    1925 => X"85",
    1926 => X"86",
    1927 => X"87",
    1928 => X"88",
    1929 => X"89",
    1930 => X"8A",
    1931 => X"8B",
    1932 => X"8C",
    1933 => X"8D",
    1934 => X"8E",
    1935 => X"8F",
    1936 => X"90",
    1937 => X"91",
    1938 => X"92",
    1939 => X"93",
    1940 => X"94",
    1941 => X"95",
    1942 => X"96",
    1943 => X"97",
    1944 => X"98",
    1945 => X"99",
    1946 => X"9A",
    1947 => X"9B",
    1948 => X"9C",
    1949 => X"9D",
    1950 => X"9E",
    1951 => X"9F",
    1952 => X"A0",
    1953 => X"A1",
    1954 => X"A2",
    1955 => X"A3",
    1956 => X"A4",
    1957 => X"A5",
    1958 => X"A6",
    1959 => X"A7",
    1960 => X"A8",
    1961 => X"A9",
    1962 => X"AA",
    1963 => X"AB",
    1964 => X"AC",
    1965 => X"AD",
    1966 => X"AE",
    1967 => X"AF",
    1968 => X"B0",
    1969 => X"B1",
    1970 => X"B2",
    1971 => X"B3",
    1972 => X"B4",
    1973 => X"B5",
    1974 => X"B6",
    1975 => X"B7",
    1976 => X"B8",
    1977 => X"B9",
    1978 => X"BA",
    1979 => X"BB",
    1980 => X"BC",
    1981 => X"BD",
    1982 => X"BE",
    1983 => X"BF",
    1984 => X"C0",
    1985 => X"C1",
    1986 => X"C2",
    1987 => X"C3",
    1988 => X"C4",
    1989 => X"C5",
    1990 => X"C6",
    1991 => X"C7",
    1992 => X"C8",
    1993 => X"C9",
    1994 => X"CA",
    1995 => X"CB",
    1996 => X"CC",
    1997 => X"CD",
    1998 => X"CE",
    1999 => X"CF",
    2000 => X"D0",
    2001 => X"D1",
    2002 => X"D2",
    2003 => X"D3",
    2004 => X"D4",
    2005 => X"D5",
    2006 => X"D6",
    2007 => X"D7",
    2008 => X"D8",
    2009 => X"D9",
    2010 => X"DA",
    2011 => X"DB",
    2012 => X"DC",
    2013 => X"DD",
    2014 => X"DE",
    2015 => X"DF",
    2016 => X"E0",
    2017 => X"E1",
    2018 => X"E2",
    2019 => X"E3",
    2020 => X"E4",
    2021 => X"E5",
    2022 => X"E6",
    2023 => X"E7",
    2024 => X"E8",
    2025 => X"E9",
    2026 => X"EA",
    2027 => X"EB",
    2028 => X"EC",
    2029 => X"ED",
    2030 => X"EE",
    2031 => X"EF",
    2032 => X"F0",
    2033 => X"F1",
    2034 => X"F2",
    2035 => X"F3",
    2036 => X"F4",
    2037 => X"F5",
    2038 => X"F6",
    2039 => X"F7",
    2040 => X"F8",
    2041 => X"F9",
    2042 => X"FA",
    2043 => X"FB",
    2044 => X"FC",
    2045 => X"FD",
    2046 => X"FE",
    2047 => X"FF",
    2048 => X"00",
    2049 => X"01",
    2050 => X"02",
    2051 => X"03",
    2052 => X"04",
    2053 => X"05",
    2054 => X"06",
    2055 => X"07",
    2056 => X"08",
    2057 => X"09",
    2058 => X"0A",
    2059 => X"0B",
    2060 => X"0C",
    2061 => X"0D",
    2062 => X"0E",
    2063 => X"0F",
    2064 => X"10",
    2065 => X"11",
    2066 => X"12",
    2067 => X"13",
    2068 => X"14",
    2069 => X"15",
    2070 => X"16",
    2071 => X"17",
    2072 => X"18",
    2073 => X"19",
    2074 => X"1A",
    2075 => X"1B",
    2076 => X"1C",
    2077 => X"1D",
    2078 => X"1E",
    2079 => X"1F",
    2080 => X"20",
    2081 => X"21",
    2082 => X"22",
    2083 => X"23",
    2084 => X"24",
    2085 => X"25",
    2086 => X"26",
    2087 => X"27",
    2088 => X"28",
    2089 => X"29",
    2090 => X"2A",
    2091 => X"2B",
    2092 => X"2C",
    2093 => X"2D",
    2094 => X"2E",
    2095 => X"2F",
    2096 => X"30",
    2097 => X"31",
    2098 => X"32",
    2099 => X"33",
    2100 => X"34",
    2101 => X"35",
    2102 => X"36",
    2103 => X"37",
    2104 => X"38",
    2105 => X"39",
    2106 => X"3A",
    2107 => X"3B",
    2108 => X"3C",
    2109 => X"3D",
    2110 => X"3E",
    2111 => X"3F",
    2112 => X"40",
    2113 => X"41",
    2114 => X"42",
    2115 => X"43",
    2116 => X"44",
    2117 => X"45",
    2118 => X"46",
    2119 => X"47",
    2120 => X"48",
    2121 => X"49",
    2122 => X"4A",
    2123 => X"4B",
    2124 => X"4C",
    2125 => X"4D",
    2126 => X"4E",
    2127 => X"4F",
    2128 => X"50",
    2129 => X"51",
    2130 => X"52",
    2131 => X"53",
    2132 => X"54",
    2133 => X"55",
    2134 => X"56",
    2135 => X"57",
    2136 => X"58",
    2137 => X"59",
    2138 => X"5A",
    2139 => X"5B",
    2140 => X"5C",
    2141 => X"5D",
    2142 => X"5E",
    2143 => X"5F",
    2144 => X"60",
    2145 => X"61",
    2146 => X"62",
    2147 => X"63",
    2148 => X"64",
    2149 => X"65",
    2150 => X"66",
    2151 => X"67",
    2152 => X"68",
    2153 => X"69",
    2154 => X"6A",
    2155 => X"6B",
    2156 => X"6C",
    2157 => X"6D",
    2158 => X"6E",
    2159 => X"6F",
    2160 => X"70",
    2161 => X"71",
    2162 => X"72",
    2163 => X"73",
    2164 => X"74",
    2165 => X"75",
    2166 => X"76",
    2167 => X"77",
    2168 => X"78",
    2169 => X"79",
    2170 => X"7A",
    2171 => X"7B",
    2172 => X"7C",
    2173 => X"7D",
    2174 => X"7E",
    2175 => X"7F",
    2176 => X"80",
    2177 => X"81",
    2178 => X"82",
    2179 => X"83",
    2180 => X"84",
    2181 => X"85",
    2182 => X"86",
    2183 => X"87",
    2184 => X"88",
    2185 => X"89",
    2186 => X"8A",
    2187 => X"8B",
    2188 => X"8C",
    2189 => X"8D",
    2190 => X"8E",
    2191 => X"8F",
    2192 => X"90",
    2193 => X"91",
    2194 => X"92",
    2195 => X"93",
    2196 => X"94",
    2197 => X"95",
    2198 => X"96",
    2199 => X"97",
    2200 => X"98",
    2201 => X"99",
    2202 => X"9A",
    2203 => X"9B",
    2204 => X"9C",
    2205 => X"9D",
    2206 => X"9E",
    2207 => X"9F",
    2208 => X"A0",
    2209 => X"A1",
    2210 => X"A2",
    2211 => X"A3",
    2212 => X"A4",
    2213 => X"A5",
    2214 => X"A6",
    2215 => X"A7",
    2216 => X"A8",
    2217 => X"A9",
    2218 => X"AA",
    2219 => X"AB",
    2220 => X"AC",
    2221 => X"AD",
    2222 => X"AE",
    2223 => X"AF",
    2224 => X"B0",
    2225 => X"B1",
    2226 => X"B2",
    2227 => X"B3",
    2228 => X"B4",
    2229 => X"B5",
    2230 => X"B6",
    2231 => X"B7",
    2232 => X"B8",
    2233 => X"B9",
    2234 => X"BA",
    2235 => X"BB",
    2236 => X"BC",
    2237 => X"BD",
    2238 => X"BE",
    2239 => X"BF",
    2240 => X"C0",
    2241 => X"C1",
    2242 => X"C2",
    2243 => X"C3",
    2244 => X"C4",
    2245 => X"C5",
    2246 => X"C6",
    2247 => X"C7",
    2248 => X"C8",
    2249 => X"C9",
    2250 => X"CA",
    2251 => X"CB",
    2252 => X"CC",
    2253 => X"CD",
    2254 => X"CE",
    2255 => X"CF",
    2256 => X"D0",
    2257 => X"D1",
    2258 => X"D2",
    2259 => X"D3",
    2260 => X"D4",
    2261 => X"D5",
    2262 => X"D6",
    2263 => X"D7",
    2264 => X"D8",
    2265 => X"D9",
    2266 => X"DA",
    2267 => X"DB",
    2268 => X"DC",
    2269 => X"DD",
    2270 => X"DE",
    2271 => X"DF",
    2272 => X"E0",
    2273 => X"E1",
    2274 => X"E2",
    2275 => X"E3",
    2276 => X"E4",
    2277 => X"E5",
    2278 => X"E6",
    2279 => X"E7",
    2280 => X"E8",
    2281 => X"E9",
    2282 => X"EA",
    2283 => X"EB",
    2284 => X"EC",
    2285 => X"ED",
    2286 => X"EE",
    2287 => X"EF",
    2288 => X"F0",
    2289 => X"F1",
    2290 => X"F2",
    2291 => X"F3",
    2292 => X"F4",
    2293 => X"F5",
    2294 => X"F6",
    2295 => X"F7",
    2296 => X"F8",
    2297 => X"F9",
    2298 => X"FA",
    2299 => X"FB",
    2300 => X"FC",
    2301 => X"FD",
    2302 => X"FE",
    2303 => X"FF",
    2304 => X"00",
    2305 => X"01",
    2306 => X"02",
    2307 => X"03",
    2308 => X"04",
    2309 => X"05",
    2310 => X"06",
    2311 => X"07",
    2312 => X"08",
    2313 => X"09",
    2314 => X"0A",
    2315 => X"0B",
    2316 => X"0C",
    2317 => X"0D",
    2318 => X"0E",
    2319 => X"0F",
    2320 => X"10",
    2321 => X"11",
    2322 => X"12",
    2323 => X"13",
    2324 => X"14",
    2325 => X"15",
    2326 => X"16",
    2327 => X"17",
    2328 => X"18",
    2329 => X"19",
    2330 => X"1A",
    2331 => X"1B",
    2332 => X"1C",
    2333 => X"1D",
    2334 => X"1E",
    2335 => X"1F",
    2336 => X"20",
    2337 => X"21",
    2338 => X"22",
    2339 => X"23",
    2340 => X"24",
    2341 => X"25",
    2342 => X"26",
    2343 => X"27",
    2344 => X"28",
    2345 => X"29",
    2346 => X"2A",
    2347 => X"2B",
    2348 => X"2C",
    2349 => X"2D",
    2350 => X"2E",
    2351 => X"2F",
    2352 => X"30",
    2353 => X"31",
    2354 => X"32",
    2355 => X"33",
    2356 => X"34",
    2357 => X"35",
    2358 => X"36",
    2359 => X"37",
    2360 => X"38",
    2361 => X"39",
    2362 => X"3A",
    2363 => X"3B",
    2364 => X"3C",
    2365 => X"3D",
    2366 => X"3E",
    2367 => X"3F",
    2368 => X"40",
    2369 => X"41",
    2370 => X"42",
    2371 => X"43",
    2372 => X"44",
    2373 => X"45",
    2374 => X"46",
    2375 => X"47",
    2376 => X"48",
    2377 => X"49",
    2378 => X"4A",
    2379 => X"4B",
    2380 => X"4C",
    2381 => X"4D",
    2382 => X"4E",
    2383 => X"4F",
    2384 => X"50",
    2385 => X"51",
    2386 => X"52",
    2387 => X"53",
    2388 => X"54",
    2389 => X"55",
    2390 => X"56",
    2391 => X"57",
    2392 => X"58",
    2393 => X"59",
    2394 => X"5A",
    2395 => X"5B",
    2396 => X"5C",
    2397 => X"5D",
    2398 => X"5E",
    2399 => X"5F",
    2400 => X"60",
    2401 => X"61",
    2402 => X"62",
    2403 => X"63",
    2404 => X"64",
    2405 => X"65",
    2406 => X"66",
    2407 => X"67",
    2408 => X"68",
    2409 => X"69",
    2410 => X"6A",
    2411 => X"6B",
    2412 => X"6C",
    2413 => X"6D",
    2414 => X"6E",
    2415 => X"6F",
    2416 => X"70",
    2417 => X"71",
    2418 => X"72",
    2419 => X"73",
    2420 => X"74",
    2421 => X"75",
    2422 => X"76",
    2423 => X"77",
    2424 => X"78",
    2425 => X"79",
    2426 => X"7A",
    2427 => X"7B",
    2428 => X"7C",
    2429 => X"7D",
    2430 => X"7E",
    2431 => X"7F",
    2432 => X"80",
    2433 => X"81",
    2434 => X"82",
    2435 => X"83",
    2436 => X"84",
    2437 => X"85",
    2438 => X"86",
    2439 => X"87",
    2440 => X"88",
    2441 => X"89",
    2442 => X"8A",
    2443 => X"8B",
    2444 => X"8C",
    2445 => X"8D",
    2446 => X"8E",
    2447 => X"8F",
    2448 => X"90",
    2449 => X"91",
    2450 => X"92",
    2451 => X"93",
    2452 => X"94",
    2453 => X"95",
    2454 => X"96",
    2455 => X"97",
    2456 => X"98",
    2457 => X"99",
    2458 => X"9A",
    2459 => X"9B",
    2460 => X"9C",
    2461 => X"9D",
    2462 => X"9E",
    2463 => X"9F",
    2464 => X"A0",
    2465 => X"A1",
    2466 => X"A2",
    2467 => X"A3",
    2468 => X"A4",
    2469 => X"A5",
    2470 => X"A6",
    2471 => X"A7",
    2472 => X"A8",
    2473 => X"A9",
    2474 => X"AA",
    2475 => X"AB",
    2476 => X"AC",
    2477 => X"AD",
    2478 => X"AE",
    2479 => X"AF",
    2480 => X"B0",
    2481 => X"B1",
    2482 => X"B2",
    2483 => X"B3",
    2484 => X"B4",
    2485 => X"B5",
    2486 => X"B6",
    2487 => X"B7",
    2488 => X"B8",
    2489 => X"B9",
    2490 => X"BA",
    2491 => X"BB",
    2492 => X"BC",
    2493 => X"BD",
    2494 => X"BE",
    2495 => X"BF",
    2496 => X"C0",
    2497 => X"C1",
    2498 => X"C2",
    2499 => X"C3",
    2500 => X"C4",
    2501 => X"C5",
    2502 => X"C6",
    2503 => X"C7",
    2504 => X"C8",
    2505 => X"C9",
    2506 => X"CA",
    2507 => X"CB",
    2508 => X"CC",
    2509 => X"CD",
    2510 => X"CE",
    2511 => X"CF",
    2512 => X"D0",
    2513 => X"D1",
    2514 => X"D2",
    2515 => X"D3",
    2516 => X"D4",
    2517 => X"D5",
    2518 => X"D6",
    2519 => X"D7",
    2520 => X"D8",
    2521 => X"D9",
    2522 => X"DA",
    2523 => X"DB",
    2524 => X"DC",
    2525 => X"DD",
    2526 => X"DE",
    2527 => X"DF",
    2528 => X"E0",
    2529 => X"E1",
    2530 => X"E2",
    2531 => X"E3",
    2532 => X"E4",
    2533 => X"E5",
    2534 => X"E6",
    2535 => X"E7",
    2536 => X"E8",
    2537 => X"E9",
    2538 => X"EA",
    2539 => X"EB",
    2540 => X"EC",
    2541 => X"ED",
    2542 => X"EE",
    2543 => X"EF",
    2544 => X"F0",
    2545 => X"F1",
    2546 => X"F2",
    2547 => X"F3",
    2548 => X"F4",
    2549 => X"F5",
    2550 => X"F6",
    2551 => X"F7",
    2552 => X"F8",
    2553 => X"F9",
    2554 => X"FA",
    2555 => X"FB",
    2556 => X"FC",
    2557 => X"FD",
    2558 => X"FE",
    2559 => X"FF",
    2560 => X"00",
    2561 => X"01",
    2562 => X"02",
    2563 => X"03",
    2564 => X"04",
    2565 => X"05",
    2566 => X"06",
    2567 => X"07",
    2568 => X"08",
    2569 => X"09",
    2570 => X"0A",
    2571 => X"0B",
    2572 => X"0C",
    2573 => X"0D",
    2574 => X"0E",
    2575 => X"0F",
    2576 => X"10",
    2577 => X"11",
    2578 => X"12",
    2579 => X"13",
    2580 => X"14",
    2581 => X"15",
    2582 => X"16",
    2583 => X"17",
    2584 => X"18",
    2585 => X"19",
    2586 => X"1A",
    2587 => X"1B",
    2588 => X"1C",
    2589 => X"1D",
    2590 => X"1E",
    2591 => X"1F",
    2592 => X"20",
    2593 => X"21",
    2594 => X"22",
    2595 => X"23",
    2596 => X"24",
    2597 => X"25",
    2598 => X"26",
    2599 => X"27",
    2600 => X"28",
    2601 => X"29",
    2602 => X"2A",
    2603 => X"2B",
    2604 => X"2C",
    2605 => X"2D",
    2606 => X"2E",
    2607 => X"2F",
    2608 => X"30",
    2609 => X"31",
    2610 => X"32",
    2611 => X"33",
    2612 => X"34",
    2613 => X"35",
    2614 => X"36",
    2615 => X"37",
    2616 => X"38",
    2617 => X"39",
    2618 => X"3A",
    2619 => X"3B",
    2620 => X"3C",
    2621 => X"3D",
    2622 => X"3E",
    2623 => X"3F",
    2624 => X"40",
    2625 => X"41",
    2626 => X"42",
    2627 => X"43",
    2628 => X"44",
    2629 => X"45",
    2630 => X"46",
    2631 => X"47",
    2632 => X"48",
    2633 => X"49",
    2634 => X"4A",
    2635 => X"4B",
    2636 => X"4C",
    2637 => X"4D",
    2638 => X"4E",
    2639 => X"4F",
    2640 => X"50",
    2641 => X"51",
    2642 => X"52",
    2643 => X"53",
    2644 => X"54",
    2645 => X"55",
    2646 => X"56",
    2647 => X"57",
    2648 => X"58",
    2649 => X"59",
    2650 => X"5A",
    2651 => X"5B",
    2652 => X"5C",
    2653 => X"5D",
    2654 => X"5E",
    2655 => X"5F",
    2656 => X"60",
    2657 => X"61",
    2658 => X"62",
    2659 => X"63",
    2660 => X"64",
    2661 => X"65",
    2662 => X"66",
    2663 => X"67",
    2664 => X"68",
    2665 => X"69",
    2666 => X"6A",
    2667 => X"6B",
    2668 => X"6C",
    2669 => X"6D",
    2670 => X"6E",
    2671 => X"6F",
    2672 => X"70",
    2673 => X"71",
    2674 => X"72",
    2675 => X"73",
    2676 => X"74",
    2677 => X"75",
    2678 => X"76",
    2679 => X"77",
    2680 => X"78",
    2681 => X"79",
    2682 => X"7A",
    2683 => X"7B",
    2684 => X"7C",
    2685 => X"7D",
    2686 => X"7E",
    2687 => X"7F",
    2688 => X"80",
    2689 => X"81",
    2690 => X"82",
    2691 => X"83",
    2692 => X"84",
    2693 => X"85",
    2694 => X"86",
    2695 => X"87",
    2696 => X"88",
    2697 => X"89",
    2698 => X"8A",
    2699 => X"8B",
    2700 => X"8C",
    2701 => X"8D",
    2702 => X"8E",
    2703 => X"8F",
    2704 => X"90",
    2705 => X"91",
    2706 => X"92",
    2707 => X"93",
    2708 => X"94",
    2709 => X"95",
    2710 => X"96",
    2711 => X"97",
    2712 => X"98",
    2713 => X"99",
    2714 => X"9A",
    2715 => X"9B",
    2716 => X"9C",
    2717 => X"9D",
    2718 => X"9E",
    2719 => X"9F",
    2720 => X"A0",
    2721 => X"A1",
    2722 => X"A2",
    2723 => X"A3",
    2724 => X"A4",
    2725 => X"A5",
    2726 => X"A6",
    2727 => X"A7",
    2728 => X"A8",
    2729 => X"A9",
    2730 => X"AA",
    2731 => X"AB",
    2732 => X"AC",
    2733 => X"AD",
    2734 => X"AE",
    2735 => X"AF",
    2736 => X"B0",
    2737 => X"B1",
    2738 => X"B2",
    2739 => X"B3",
    2740 => X"B4",
    2741 => X"B5",
    2742 => X"B6",
    2743 => X"B7",
    2744 => X"B8",
    2745 => X"B9",
    2746 => X"BA",
    2747 => X"BB",
    2748 => X"BC",
    2749 => X"BD",
    2750 => X"BE",
    2751 => X"BF",
    2752 => X"C0",
    2753 => X"C1",
    2754 => X"C2",
    2755 => X"C3",
    2756 => X"C4",
    2757 => X"C5",
    2758 => X"C6",
    2759 => X"C7",
    2760 => X"C8",
    2761 => X"C9",
    2762 => X"CA",
    2763 => X"CB",
    2764 => X"CC",
    2765 => X"CD",
    2766 => X"CE",
    2767 => X"CF",
    2768 => X"D0",
    2769 => X"D1",
    2770 => X"D2",
    2771 => X"D3",
    2772 => X"D4",
    2773 => X"D5",
    2774 => X"D6",
    2775 => X"D7",
    2776 => X"D8",
    2777 => X"D9",
    2778 => X"DA",
    2779 => X"DB",
    2780 => X"DC",
    2781 => X"DD",
    2782 => X"DE",
    2783 => X"DF",
    2784 => X"E0",
    2785 => X"E1",
    2786 => X"E2",
    2787 => X"E3",
    2788 => X"E4",
    2789 => X"E5",
    2790 => X"E6",
    2791 => X"E7",
    2792 => X"E8",
    2793 => X"E9",
    2794 => X"EA",
    2795 => X"EB",
    2796 => X"EC",
    2797 => X"ED",
    2798 => X"EE",
    2799 => X"EF",
    2800 => X"F0",
    2801 => X"F1",
    2802 => X"F2",
    2803 => X"F3",
    2804 => X"F4",
    2805 => X"F5",
    2806 => X"F6",
    2807 => X"F7",
    2808 => X"F8",
    2809 => X"F9",
    2810 => X"FA",
    2811 => X"FB",
    2812 => X"FC",
    2813 => X"FD",
    2814 => X"FE",
    2815 => X"FF",
    2816 => X"00",
    2817 => X"01",
    2818 => X"02",
    2819 => X"03",
    2820 => X"04",
    2821 => X"05",
    2822 => X"06",
    2823 => X"07",
    2824 => X"08",
    2825 => X"09",
    2826 => X"0A",
    2827 => X"0B",
    2828 => X"0C",
    2829 => X"0D",
    2830 => X"0E",
    2831 => X"0F",
    2832 => X"10",
    2833 => X"11",
    2834 => X"12",
    2835 => X"13",
    2836 => X"14",
    2837 => X"15",
    2838 => X"16",
    2839 => X"17",
    2840 => X"18",
    2841 => X"19",
    2842 => X"1A",
    2843 => X"1B",
    2844 => X"1C",
    2845 => X"1D",
    2846 => X"1E",
    2847 => X"1F",
    2848 => X"20",
    2849 => X"21",
    2850 => X"22",
    2851 => X"23",
    2852 => X"24",
    2853 => X"25",
    2854 => X"26",
    2855 => X"27",
    2856 => X"28",
    2857 => X"29",
    2858 => X"2A",
    2859 => X"2B",
    2860 => X"2C",
    2861 => X"2D",
    2862 => X"2E",
    2863 => X"2F",
    2864 => X"30",
    2865 => X"31",
    2866 => X"32",
    2867 => X"33",
    2868 => X"34",
    2869 => X"35",
    2870 => X"36",
    2871 => X"37",
    2872 => X"38",
    2873 => X"39",
    2874 => X"3A",
    2875 => X"3B",
    2876 => X"3C",
    2877 => X"3D",
    2878 => X"3E",
    2879 => X"3F",
    2880 => X"40",
    2881 => X"41",
    2882 => X"42",
    2883 => X"43",
    2884 => X"44",
    2885 => X"45",
    2886 => X"46",
    2887 => X"47",
    2888 => X"48",
    2889 => X"49",
    2890 => X"4A",
    2891 => X"4B",
    2892 => X"4C",
    2893 => X"4D",
    2894 => X"4E",
    2895 => X"4F",
    2896 => X"50",
    2897 => X"51",
    2898 => X"52",
    2899 => X"53",
    2900 => X"54",
    2901 => X"55",
    2902 => X"56",
    2903 => X"57",
    2904 => X"58",
    2905 => X"59",
    2906 => X"5A",
    2907 => X"5B",
    2908 => X"5C",
    2909 => X"5D",
    2910 => X"5E",
    2911 => X"5F",
    2912 => X"60",
    2913 => X"61",
    2914 => X"62",
    2915 => X"63",
    2916 => X"64",
    2917 => X"65",
    2918 => X"66",
    2919 => X"67",
    2920 => X"68",
    2921 => X"69",
    2922 => X"6A",
    2923 => X"6B",
    2924 => X"6C",
    2925 => X"6D",
    2926 => X"6E",
    2927 => X"6F",
    2928 => X"70",
    2929 => X"71",
    2930 => X"72",
    2931 => X"73",
    2932 => X"74",
    2933 => X"75",
    2934 => X"76",
    2935 => X"77",
    2936 => X"78",
    2937 => X"79",
    2938 => X"7A",
    2939 => X"7B",
    2940 => X"7C",
    2941 => X"7D",
    2942 => X"7E",
    2943 => X"7F",
    2944 => X"80",
    2945 => X"81",
    2946 => X"82",
    2947 => X"83",
    2948 => X"84",
    2949 => X"85",
    2950 => X"86",
    2951 => X"87",
    2952 => X"88",
    2953 => X"89",
    2954 => X"8A",
    2955 => X"8B",
    2956 => X"8C",
    2957 => X"8D",
    2958 => X"8E",
    2959 => X"8F",
    2960 => X"90",
    2961 => X"91",
    2962 => X"92",
    2963 => X"93",
    2964 => X"94",
    2965 => X"95",
    2966 => X"96",
    2967 => X"97",
    2968 => X"98",
    2969 => X"99",
    2970 => X"9A",
    2971 => X"9B",
    2972 => X"9C",
    2973 => X"9D",
    2974 => X"9E",
    2975 => X"9F",
    2976 => X"A0",
    2977 => X"A1",
    2978 => X"A2",
    2979 => X"A3",
    2980 => X"A4",
    2981 => X"A5",
    2982 => X"A6",
    2983 => X"A7",
    2984 => X"A8",
    2985 => X"A9",
    2986 => X"AA",
    2987 => X"AB",
    2988 => X"AC",
    2989 => X"AD",
    2990 => X"AE",
    2991 => X"AF",
    2992 => X"B0",
    2993 => X"B1",
    2994 => X"B2",
    2995 => X"B3",
    2996 => X"B4",
    2997 => X"B5",
    2998 => X"B6",
    2999 => X"B7",
    3000 => X"B8",
    3001 => X"B9",
    3002 => X"BA",
    3003 => X"BB",
    3004 => X"BC",
    3005 => X"BD",
    3006 => X"BE",
    3007 => X"BF",
    3008 => X"C0",
    3009 => X"C1",
    3010 => X"C2",
    3011 => X"C3",
    3012 => X"C4",
    3013 => X"C5",
    3014 => X"C6",
    3015 => X"C7",
    3016 => X"C8",
    3017 => X"C9",
    3018 => X"CA",
    3019 => X"CB",
    3020 => X"CC",
    3021 => X"CD",
    3022 => X"CE",
    3023 => X"CF",
    3024 => X"D0",
    3025 => X"D1",
    3026 => X"D2",
    3027 => X"D3",
    3028 => X"D4",
    3029 => X"D5",
    3030 => X"D6",
    3031 => X"D7",
    3032 => X"D8",
    3033 => X"D9",
    3034 => X"DA",
    3035 => X"DB",
    3036 => X"DC",
    3037 => X"DD",
    3038 => X"DE",
    3039 => X"DF",
    3040 => X"E0",
    3041 => X"E1",
    3042 => X"E2",
    3043 => X"E3",
    3044 => X"E4",
    3045 => X"E5",
    3046 => X"E6",
    3047 => X"E7",
    3048 => X"E8",
    3049 => X"E9",
    3050 => X"EA",
    3051 => X"EB",
    3052 => X"EC",
    3053 => X"ED",
    3054 => X"EE",
    3055 => X"EF",
    3056 => X"F0",
    3057 => X"F1",
    3058 => X"F2",
    3059 => X"F3",
    3060 => X"F4",
    3061 => X"F5",
    3062 => X"F6",
    3063 => X"F7",
    3064 => X"F8",
    3065 => X"F9",
    3066 => X"FA",
    3067 => X"FB",
    3068 => X"FC",
    3069 => X"FD",
    3070 => X"FE",
    3071 => X"FF",
    others => (others => '0'));
end ROM_Package;